`timescale 1ns / 1ps

module Shift_reg(
    input rst,
    input clk,          // Work at 100MHz clock

    input [31:0] din,   // Data input  
    input [3:0] hex,    // Hexadecimal code for the switches
    input add,          // Add signal
    input del,          // Delete signal
    input set,          // Set signal
    
    output reg [31:0] dout  // Data output
);
//wire add1,del1;
    // TODO
//dedge_signal de(.clk(clk),.in(add),.out(add1));
//dedge_signal de1(.clk(clk),.in(del),.out(del1));
always @(posedge clk or posedge rst)
begin
if(rst)
dout <= 0;
else if(set)
dout<=din;
else
    begin
        if(add)
            dout<=(dout<<4)+hex;
        else if(del)
            dout<=(dout>>4);
    end
end
endmodule

